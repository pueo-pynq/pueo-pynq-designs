module Gaussian12b_LFSR #(parameter SEED_BASE=0)
    (
    input clk,
    input rst_i,
    output [127:0] sim_data
    );

    reg [7:0][11:0] gauss_idx;
    // wire [7:0][5:0] linear_section;
    reg [4097:0][11:0] gaussian_lut = {12'b111101101010, 12'b111101110010, 12'b111101111001, 12'b111101111110, 12'b111110000010, 12'b111110000100, 12'b111110000111, 12'b111110001001, 12'b111110001010, 12'b111110001100, 12'b111110001101, 12'b111110001110, 12'b111110010000, 12'b111110010001, 12'b111110010010, 12'b111110010011, 12'b111110010100, 12'b111110010100, 12'b111110010101, 12'b111110010110, 12'b111110010111, 12'b111110010111, 12'b111110011000, 12'b111110011001, 12'b111110011001, 12'b111110011010, 12'b111110011010, 12'b111110011011, 12'b111110011100, 12'b111110011100, 12'b111110011101, 12'b111110011101, 12'b111110011110, 12'b111110011110, 12'b111110011110, 12'b111110011111, 12'b111110011111, 12'b111110100000, 12'b111110100000, 12'b111110100000, 12'b111110100001, 12'b111110100001, 12'b111110100010, 12'b111110100010, 12'b111110100010, 12'b111110100011, 12'b111110100011, 12'b111110100011, 12'b111110100100, 12'b111110100100, 12'b111110100100, 12'b111110100101, 12'b111110100101, 12'b111110100101, 12'b111110100110, 12'b111110100110, 12'b111110100110, 12'b111110100110, 12'b111110100111, 12'b111110100111, 12'b111110100111, 12'b111110101000, 12'b111110101000, 12'b111110101000, 12'b111110101000, 12'b111110101001, 12'b111110101001, 12'b111110101001, 12'b111110101001, 12'b111110101010, 12'b111110101010, 12'b111110101010, 12'b111110101010, 12'b111110101010, 12'b111110101011, 12'b111110101011, 12'b111110101011, 12'b111110101011, 12'b111110101100, 12'b111110101100, 12'b111110101100, 12'b111110101100, 12'b111110101100, 12'b111110101101, 12'b111110101101, 12'b111110101101, 12'b111110101101, 12'b111110101101, 12'b111110101110, 12'b111110101110, 12'b111110101110, 12'b111110101110, 12'b111110101110, 12'b111110101111, 12'b111110101111, 12'b111110101111, 12'b111110101111, 12'b111110101111, 12'b111110101111, 12'b111110110000, 12'b111110110000, 12'b111110110000, 12'b111110110000, 12'b111110110000, 12'b111110110001, 12'b111110110001, 12'b111110110001, 12'b111110110001, 12'b111110110001, 12'b111110110001, 12'b111110110010, 12'b111110110010, 12'b111110110010, 12'b111110110010, 12'b111110110010, 12'b111110110010, 12'b111110110010, 12'b111110110011, 12'b111110110011, 12'b111110110011, 12'b111110110011, 12'b111110110011, 12'b111110110011, 12'b111110110011, 12'b111110110100, 12'b111110110100, 12'b111110110100, 12'b111110110100, 12'b111110110100, 12'b111110110100, 12'b111110110101, 12'b111110110101, 12'b111110110101, 12'b111110110101, 12'b111110110101, 12'b111110110101, 12'b111110110101, 12'b111110110101, 12'b111110110110, 12'b111110110110, 12'b111110110110, 12'b111110110110, 12'b111110110110, 12'b111110110110, 12'b111110110110, 12'b111110110111, 12'b111110110111, 12'b111110110111, 12'b111110110111, 12'b111110110111, 12'b111110110111, 12'b111110110111, 12'b111110110111, 12'b111110111000, 12'b111110111000, 12'b111110111000, 12'b111110111000, 12'b111110111000, 12'b111110111000, 12'b111110111000, 12'b111110111000, 12'b111110111000, 12'b111110111001, 12'b111110111001, 12'b111110111001, 12'b111110111001, 12'b111110111001, 12'b111110111001, 12'b111110111001, 12'b111110111001, 12'b111110111010, 12'b111110111010, 12'b111110111010, 12'b111110111010, 12'b111110111010, 12'b111110111010, 12'b111110111010, 12'b111110111010, 12'b111110111010, 12'b111110111011, 12'b111110111011, 12'b111110111011, 12'b111110111011, 12'b111110111011, 12'b111110111011, 12'b111110111011, 12'b111110111011, 12'b111110111011, 12'b111110111011, 12'b111110111100, 12'b111110111100, 12'b111110111100, 12'b111110111100, 12'b111110111100, 12'b111110111100, 12'b111110111100, 12'b111110111100, 12'b111110111100, 12'b111110111100, 12'b111110111101, 12'b111110111101, 12'b111110111101, 12'b111110111101, 12'b111110111101, 12'b111110111101, 12'b111110111101, 12'b111110111101, 12'b111110111101, 12'b111110111101, 12'b111110111110, 12'b111110111110, 12'b111110111110, 12'b111110111110, 12'b111110111110, 12'b111110111110, 12'b111110111110, 12'b111110111110, 12'b111110111110, 12'b111110111110, 12'b111110111110, 12'b111110111111, 12'b111110111111, 12'b111110111111, 12'b111110111111, 12'b111110111111, 12'b111110111111, 12'b111110111111, 12'b111110111111, 12'b111110111111, 12'b111110111111, 12'b111110111111, 12'b111111000000, 12'b111111000000, 12'b111111000000, 12'b111111000000, 12'b111111000000, 12'b111111000000, 12'b111111000000, 12'b111111000000, 12'b111111000000, 12'b111111000000, 12'b111111000000, 12'b111111000001, 12'b111111000001, 12'b111111000001, 12'b111111000001, 12'b111111000001, 12'b111111000001, 12'b111111000001, 12'b111111000001, 12'b111111000001, 12'b111111000001, 12'b111111000001, 12'b111111000001, 12'b111111000010, 12'b111111000010, 12'b111111000010, 12'b111111000010, 12'b111111000010, 12'b111111000010, 12'b111111000010, 12'b111111000010, 12'b111111000010, 12'b111111000010, 12'b111111000010, 12'b111111000010, 12'b111111000010, 12'b111111000011, 12'b111111000011, 12'b111111000011, 12'b111111000011, 12'b111111000011, 12'b111111000011, 12'b111111000011, 12'b111111000011, 12'b111111000011, 12'b111111000011, 12'b111111000011, 12'b111111000011, 12'b111111000011, 12'b111111000100, 12'b111111000100, 12'b111111000100, 12'b111111000100, 12'b111111000100, 12'b111111000100, 12'b111111000100, 12'b111111000100, 12'b111111000100, 12'b111111000100, 12'b111111000100, 12'b111111000100, 12'b111111000100, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000101, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000110, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111000111, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001000, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001001, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001010, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001011, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001100, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001101, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001110, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111001111, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010000, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010001, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010010, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010011, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010100, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010101, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010110, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111010111, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011000, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011001, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011010, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011011, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011100, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011101, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011110, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111011111, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100001, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100010, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100011, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100100, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100101, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100110, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111100111, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101000, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101001, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101010, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101011, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101100, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101101, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101110, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111101111, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110001, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110010, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110011, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110100, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110101, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110110, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111110111, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111000, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111001, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111010, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111011, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111100, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111101, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111110, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b111111111111, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000001, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000010, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000011, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000100, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000101, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000110, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000000111, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001000, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001001, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001010, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001011, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001100, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001101, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001110, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000001111, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010001, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010010, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010011, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010100, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010101, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010110, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000010111, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011000, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011001, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011010, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011011, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011100, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011101, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011110, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000011111, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100001, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100010, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100011, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100100, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100101, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100110, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000100111, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101000, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101001, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101010, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101011, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101100, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101101, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101110, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000101111, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110000, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110001, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110010, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110011, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110100, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110101, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110110, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000110111, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111000, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111001, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111010, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111011, 12'b000000111100, 12'b000000111100, 12'b000000111100, 12'b000000111100, 12'b000000111100, 12'b000000111100, 12'b000000111100, 12'b000000111100, 12'b000000111100, 12'b000000111100, 12'b000000111100, 12'b000000111100, 12'b000000111100, 12'b000000111101, 12'b000000111101, 12'b000000111101, 12'b000000111101, 12'b000000111101, 12'b000000111101, 12'b000000111101, 12'b000000111101, 12'b000000111101, 12'b000000111101, 12'b000000111101, 12'b000000111101, 12'b000000111101, 12'b000000111110, 12'b000000111110, 12'b000000111110, 12'b000000111110, 12'b000000111110, 12'b000000111110, 12'b000000111110, 12'b000000111110, 12'b000000111110, 12'b000000111110, 12'b000000111110, 12'b000000111110, 12'b000000111110, 12'b000000111111, 12'b000000111111, 12'b000000111111, 12'b000000111111, 12'b000000111111, 12'b000000111111, 12'b000000111111, 12'b000000111111, 12'b000000111111, 12'b000000111111, 12'b000000111111, 12'b000000111111, 12'b000001000000, 12'b000001000000, 12'b000001000000, 12'b000001000000, 12'b000001000000, 12'b000001000000, 12'b000001000000, 12'b000001000000, 12'b000001000000, 12'b000001000000, 12'b000001000000, 12'b000001000001, 12'b000001000001, 12'b000001000001, 12'b000001000001, 12'b000001000001, 12'b000001000001, 12'b000001000001, 12'b000001000001, 12'b000001000001, 12'b000001000001, 12'b000001000001, 12'b000001000010, 12'b000001000010, 12'b000001000010, 12'b000001000010, 12'b000001000010, 12'b000001000010, 12'b000001000010, 12'b000001000010, 12'b000001000010, 12'b000001000010, 12'b000001000010, 12'b000001000011, 12'b000001000011, 12'b000001000011, 12'b000001000011, 12'b000001000011, 12'b000001000011, 12'b000001000011, 12'b000001000011, 12'b000001000011, 12'b000001000011, 12'b000001000100, 12'b000001000100, 12'b000001000100, 12'b000001000100, 12'b000001000100, 12'b000001000100, 12'b000001000100, 12'b000001000100, 12'b000001000100, 12'b000001000100, 12'b000001000101, 12'b000001000101, 12'b000001000101, 12'b000001000101, 12'b000001000101, 12'b000001000101, 12'b000001000101, 12'b000001000101, 12'b000001000101, 12'b000001000101, 12'b000001000110, 12'b000001000110, 12'b000001000110, 12'b000001000110, 12'b000001000110, 12'b000001000110, 12'b000001000110, 12'b000001000110, 12'b000001000110, 12'b000001000111, 12'b000001000111, 12'b000001000111, 12'b000001000111, 12'b000001000111, 12'b000001000111, 12'b000001000111, 12'b000001000111, 12'b000001001000, 12'b000001001000, 12'b000001001000, 12'b000001001000, 12'b000001001000, 12'b000001001000, 12'b000001001000, 12'b000001001000, 12'b000001001000, 12'b000001001001, 12'b000001001001, 12'b000001001001, 12'b000001001001, 12'b000001001001, 12'b000001001001, 12'b000001001001, 12'b000001001001, 12'b000001001010, 12'b000001001010, 12'b000001001010, 12'b000001001010, 12'b000001001010, 12'b000001001010, 12'b000001001010, 12'b000001001011, 12'b000001001011, 12'b000001001011, 12'b000001001011, 12'b000001001011, 12'b000001001011, 12'b000001001011, 12'b000001001011, 12'b000001001100, 12'b000001001100, 12'b000001001100, 12'b000001001100, 12'b000001001100, 12'b000001001100, 12'b000001001101, 12'b000001001101, 12'b000001001101, 12'b000001001101, 12'b000001001101, 12'b000001001101, 12'b000001001101, 12'b000001001110, 12'b000001001110, 12'b000001001110, 12'b000001001110, 12'b000001001110, 12'b000001001110, 12'b000001001110, 12'b000001001111, 12'b000001001111, 12'b000001001111, 12'b000001001111, 12'b000001001111, 12'b000001001111, 12'b000001010000, 12'b000001010000, 12'b000001010000, 12'b000001010000, 12'b000001010000, 12'b000001010001, 12'b000001010001, 12'b000001010001, 12'b000001010001, 12'b000001010001, 12'b000001010001, 12'b000001010010, 12'b000001010010, 12'b000001010010, 12'b000001010010, 12'b000001010010, 12'b000001010011, 12'b000001010011, 12'b000001010011, 12'b000001010011, 12'b000001010011, 12'b000001010100, 12'b000001010100, 12'b000001010100, 12'b000001010100, 12'b000001010100, 12'b000001010101, 12'b000001010101, 12'b000001010101, 12'b000001010101, 12'b000001010110, 12'b000001010110, 12'b000001010110, 12'b000001010110, 12'b000001010110, 12'b000001010111, 12'b000001010111, 12'b000001010111, 12'b000001010111, 12'b000001011000, 12'b000001011000, 12'b000001011000, 12'b000001011000, 12'b000001011001, 12'b000001011001, 12'b000001011001, 12'b000001011010, 12'b000001011010, 12'b000001011010, 12'b000001011010, 12'b000001011011, 12'b000001011011, 12'b000001011011, 12'b000001011100, 12'b000001011100, 12'b000001011100, 12'b000001011101, 12'b000001011101, 12'b000001011101, 12'b000001011110, 12'b000001011110, 12'b000001011110, 12'b000001011111, 12'b000001011111, 12'b000001100000, 12'b000001100000, 12'b000001100000, 12'b000001100001, 12'b000001100001, 12'b000001100010, 12'b000001100010, 12'b000001100010, 12'b000001100011, 12'b000001100011, 12'b000001100100, 12'b000001100100, 12'b000001100101, 12'b000001100110, 12'b000001100110, 12'b000001100111, 12'b000001100111, 12'b000001101000, 12'b000001101001, 12'b000001101001, 12'b000001101010, 12'b000001101011, 12'b000001101100, 12'b000001101100, 12'b000001101101, 12'b000001101110, 12'b000001101111, 12'b000001110000, 12'b000001110010, 12'b000001110011, 12'b000001110100, 12'b000001110110, 12'b000001110111, 12'b000001111001, 12'b000001111100, 12'b000001111110, 12'b000010000010, 12'b000010000111, 12'b000010001110};

    genvar idx;
    generate
        for(idx=0; idx<8; idx++) begin
            LFSR #(.NUM_BITS(12)) LFSR_idx( .i_Clk(clk),
                                            .i_Enable(1'b1),
                                            .i_Seed_DV(rst_i),
                                            .i_Seed_Data(SEED_BASE+idx*256),
                                            .o_LFSR_Data(gauss_idx[idx])
                                            );


            assign sim_data[(idx*16) +: 12]      = gaussian_lut[gauss_idx[idx]];
            assign sim_data[(idx*16 + 12) +: 4] = {4{gaussian_lut[gauss_idx[idx]][11]}};
        end
    endgenerate
    

endmodule