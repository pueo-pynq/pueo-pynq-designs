module Gaussian12b_LFSR #(parameter SEED_BASE=0)
    (
    input clk,
    output [127:0] sim_data
    );

    reg [7:0][7:0] gauss_idx;
    wire [7:0][5:0] linear_section;
    reg [255:0][11:0] gaussian_lut = {12'b100100010000, 12'b100110110000, 12'b101001000000, 12'b101010100000, 12'b101011100000, 12'b101100100000, 12'b101101000000, 12'b101101110000, 12'b101110010000, 12'b101110110000, 12'b101111010000, 12'b101111110000, 12'b110000000000, 12'b110000100000, 12'b110000110000, 12'b110001010000, 12'b110001100000, 12'b110001110000, 12'b110010000000, 12'b110010010000, 12'b110010100000, 12'b110010110000, 12'b110011000000, 12'b110011010000, 12'b110011100000, 12'b110011110000, 12'b110100000000, 12'b110100010000, 12'b110100010000, 12'b110100100000, 12'b110100110000, 12'b110101000000, 12'b110101000000, 12'b110101010000, 12'b110101100000, 12'b110101110000, 12'b110101110000, 12'b110110000000, 12'b110110010000, 12'b110110010000, 12'b110110100000, 12'b110110100000, 12'b110110110000, 12'b110111000000, 12'b110111000000, 12'b110111010000, 12'b110111010000, 12'b110111100000, 12'b110111110000, 12'b110111110000, 12'b111000000000, 12'b111000000000, 12'b111000010000, 12'b111000010000, 12'b111000100000, 12'b111000100000, 12'b111000110000, 12'b111000110000, 12'b111001000000, 12'b111001000000, 12'b111001010000, 12'b111001010000, 12'b111001100000, 12'b111001100000, 12'b111001110000, 12'b111001110000, 12'b111010000000, 12'b111010000000, 12'b111010010000, 12'b111010010000, 12'b111010010000, 12'b111010100000, 12'b111010100000, 12'b111010110000, 12'b111010110000, 12'b111011000000, 12'b111011000000, 12'b111011010000, 12'b111011010000, 12'b111011010000, 12'b111011100000, 12'b111011100000, 12'b111011110000, 12'b111011110000, 12'b111011110000, 12'b111100000000, 12'b111100000000, 12'b111100010000, 12'b111100010000, 12'b111100100000, 12'b111100100000, 12'b111100100000, 12'b111100110000, 12'b111100110000, 12'b111101000000, 12'b111101000000, 12'b111101000000, 12'b111101010000, 12'b111101010000, 12'b111101010000, 12'b111101100000, 12'b111101100000, 12'b111101110000, 12'b111101110000, 12'b111101110000, 12'b111110000000, 12'b111110000000, 12'b111110010000, 12'b111110010000, 12'b111110010000, 12'b111110100000, 12'b111110100000, 12'b111110100000, 12'b111110110000, 12'b111110110000, 12'b111111000000, 12'b111111000000, 12'b111111000000, 12'b111111010000, 12'b111111010000, 12'b111111100000, 12'b111111100000, 12'b111111100000, 12'b111111110000, 12'b111111110000, 12'b111111110000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000000000, 12'b000000010000, 12'b000000010000, 12'b000000010000, 12'b000000100000, 12'b000000100000, 12'b000000100000, 12'b000000110000, 12'b000000110000, 12'b000001000000, 12'b000001000000, 12'b000001000000, 12'b000001010000, 12'b000001010000, 12'b000001100000, 12'b000001100000, 12'b000001100000, 12'b000001110000, 12'b000001110000, 12'b000001110000, 12'b000010000000, 12'b000010000000, 12'b000010010000, 12'b000010010000, 12'b000010010000, 12'b000010100000, 12'b000010100000, 12'b000010110000, 12'b000010110000, 12'b000010110000, 12'b000011000000, 12'b000011000000, 12'b000011000000, 12'b000011010000, 12'b000011010000, 12'b000011100000, 12'b000011100000, 12'b000011100000, 12'b000011110000, 12'b000011110000, 12'b000100000000, 12'b000100000000, 12'b000100010000, 12'b000100010000, 12'b000100010000, 12'b000100100000, 12'b000100100000, 12'b000100110000, 12'b000100110000, 12'b000100110000, 12'b000101000000, 12'b000101000000, 12'b000101010000, 12'b000101010000, 12'b000101100000, 12'b000101100000, 12'b000101110000, 12'b000101110000, 12'b000101110000, 12'b000110000000, 12'b000110000000, 12'b000110010000, 12'b000110010000, 12'b000110100000, 12'b000110100000, 12'b000110110000, 12'b000110110000, 12'b000111000000, 12'b000111000000, 12'b000111010000, 12'b000111010000, 12'b000111100000, 12'b000111100000, 12'b000111110000, 12'b000111110000, 12'b001000000000, 12'b001000000000, 12'b001000010000, 12'b001000010000, 12'b001000100000, 12'b001000110000, 12'b001000110000, 12'b001001000000, 12'b001001000000, 12'b001001010000, 12'b001001100000, 12'b001001100000, 12'b001001110000, 12'b001001110000, 12'b001010000000, 12'b001010010000, 12'b001010010000, 12'b001010100000, 12'b001010110000, 12'b001011000000, 12'b001011000000, 12'b001011010000, 12'b001011100000, 12'b001011110000, 12'b001011110000, 12'b001100000000, 12'b001100010000, 12'b001100100000, 12'b001100110000, 12'b001101000000, 12'b001101010000, 12'b001101100000, 12'b001101110000, 12'b001110000000, 12'b001110010000, 12'b001110100000, 12'b001110110000, 12'b001111010000, 12'b001111100000, 12'b010000000000, 12'b010000010000, 12'b010000110000, 12'b010001010000, 12'b010001110000, 12'b010010010000, 12'b010011000000, 12'b010011100000, 12'b010100100000, 12'b010101100000, 12'b010111000000, 12'b011001010000};

    genvar idx;
    generate
        for(idx=0; idx<8; idx++) begin
            LFSR #(.NUM_BITS(8)) LFSR_idx( .i_Clk(clk),
                                            .i_Enable(1'b1),
                                            .i_Seed_DV(1'b0),
                                            .i_Seed_Data(SEED_BASE+idx+1),
                                            .o_LFSR_Data(gauss_idx[idx])
                                            );

            LFSR #(.NUM_BITS(6)) LFSR_lin( .i_Clk(clk),
                                            .i_Enable(1'b1),
                                            .i_Seed_DV(1'b1),
                                            .i_Seed_Data(SEED_BASE+idx+16),
                                            .o_LFSR_Data(linear_section[idx])
                                            );

            
            // assign sim_data[(idx*16 + 8) +: 8]    = gaussian_lut[gauss_idx][4+:8];
            // assign sim_data[(idx*16 + 4) +: 4]    = linear_section[idx];
            // assign sim_data[idx*16 +: 4]          = 4'b0000;
            assign sim_data[(idx*16) +: 6]      = linear_section[gauss_idx][5:0];
            assign sim_data[(idx*16+6) +: 8]    = gaussian_lut[gauss_idx][4+:8];
            assign sim_data[(idx*16 + 14) +: 2] = {2{gaussian_lut[gauss_idx][11]}};
        end
    endgenerate
    

endmodule